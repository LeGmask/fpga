-- fichier à écraser avec le fichier de test généré par ISE (New Source)
-- le nom du composant de test doit être TestOpl (respect minuscules/majuscules)
