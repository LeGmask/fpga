../er_1octet/er_1octet.vhd